
module IVS_ONEHOT_BIN_SEL(/*autoarg*/
    // Outputs
    bin,
    // Inputs
    ori
    );
    input [31:0]    ori;
    output [ 31:0]  bin;

    assign bin = ori[ 0] ? 32'h0000_0001 :
                 ori[ 1] ? 32'h0000_0002 :
                 ori[ 2] ? 32'h0000_0004 :
                 ori[ 3] ? 32'h0000_0008 :
                 ori[ 4] ? 32'h0000_0010 :
                 ori[ 5] ? 32'h0000_0020 :
                 ori[ 6] ? 32'h0000_0040 :
                 ori[ 7] ? 32'h0000_0080 :
                 ori[ 8] ? 32'h0000_0100 :
                 ori[ 9] ? 32'h0000_0200 :
                 ori[10] ? 32'h0000_0400 :
                 ori[11] ? 32'h0000_0800 :
                 ori[12] ? 32'h0000_1000 :
                 ori[13] ? 32'h0000_2000 :
                 ori[14] ? 32'h0000_4000 :
                 ori[15] ? 32'h0000_8000 :
                 ori[16] ? 32'h0001_0000 :
                 ori[17] ? 32'h0002_0000 :
                 ori[18] ? 32'h0004_0000 :
                 ori[19] ? 32'h0008_0000 :
                 ori[20] ? 32'h0010_0000 :
                 ori[21] ? 32'h0020_0000 :
                 ori[22] ? 32'h0040_0000 :
                 ori[23] ? 32'h0080_0000 :
                 ori[24] ? 32'h0100_0000 :
                 ori[25] ? 32'h0200_0000 :
                 ori[26] ? 32'h0400_0000 :
                 ori[27] ? 32'h0800_0000 :
                 ori[28] ? 32'h1000_0000 :
                 ori[29] ? 32'h2000_0000 :
                 ori[30] ? 32'h4000_0000 :
                 ori[31] ? 32'h8000_0000 : 32'h0000_0000;
    
    
endmodule // IVS_ONEHOT_BIN_SEL

